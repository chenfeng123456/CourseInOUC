LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY homework3 IS
   PORT ( 
	       clk, dir: IN STD_LOGIC;
	       a, b, c, d: OUT STD_LOGIC
		  );
END;

ARCHITECTURE bhv OF homework3 IS
BEGIN
END;